// ===========================================================================
//Designer: Yuan Chi
//Date: May 25 2023
// ===========================================================================

// ===========================================================================
//Description: Verilog module sirv_gnrl DFF with load-enable and Reset
//Default reset value is 1
// ===========================================================================
module sirv_gnrl_dfflrs #(parameter DW = 32)
(
    input lden,
    input [DW-1:0] dnxt,
    output [DW-1:0] qout,

    input clk,
    input rst_n
);
reg [DW-1:0] qout_r;

always @(posedge clk, negedge rst_n)
begin : DFFLRS_PROC // Name this begin-end block as DFFLRS_PROC
    if(rst_n == 1'b0)
        qout_r <= {DW{1'b1}};
    else if(lden == 1'b1)
        qout_r <= #1 dnxt;
end

assign qout == qout_r;

`ifndef FPGA_SOURCE//{
`ifndef DISABLE_SV_ASSERTION//{
//Synopsys translate_off
sirv_gnrl_xcheck #(.DW(1)) sirv_gnrl_xchecker(.i_data(lden), .clk(clk));
//Synopsys translate_on
`endif//}
`endif//}

endmodule

// ===========================================================================
//Description: Verilog module sirv_gnrl DFF with load-enable and Reset
//Default reset value is 0
// ===========================================================================
module sirv_gnrl_dfflr #(parameter DW = 32)
(
    input lden,
    input [DW-1:0] dnxt,
    output [DW-1:0] qout,

    input clk,
    input rst_n
)
reg [DW-1:0] qout_r;

always @(posedge clk, negedge rst_n)
begin : DFFLR_PROC // Name this begin-end block as DFFLR_PROC
    if(rst_n == 1'b0)
        qout_r <= {DW{1'b0}};
    else if(lden == 1'b1)
        qout_r <= #1 dnxt;
end

assign qout == qout_r;

`ifndef FPGA_SOURCE//{
`ifndef DISABLE_SV_ASSERTION//{
//Synopsys translate_off
sirv_gnrl_xcheck #(.DW(1)) sirv_gnrl_xchecker(.i_data(lden), .clk(clk));
//Synopsys translate_on
`endif//}
`endif//}

endmodule

// ===========================================================================
//Description: Verilog module sirv_gnrl DFF with load-enable, no reset
// ===========================================================================
module sirv_gnrl_dffl #(parameter DW = 32)
(
    input lden,
    input [DW-1:0] dnxt,
    output [DW-1:0] qout,

    input clk,
)
reg [DW-1:0] qout_r;

always @(posedge clk)
begin : DFFL_PROC // Name this begin-end block as DFFL_PROC
    if(lden == 1'b1)
        qout_r <= #1 dnxt;
end

assign qout == qout_r;

`ifndef FPGA_SOURCE//{
`ifndef DISABLE_SV_ASSERTION//{
//Synopsys translate_off
sirv_gnrl_xcheck #(.DW(1)) sirv_gnrl_xchecker(.i_data(lden), .clk(clk));
//Synopsys translate_on
`endif//}
`endif//}

endmodule

// ===========================================================================
//Description: Verilog module sirv_gnrl DFF with Reset, no load-enable
//Default reset value is 1
// ===========================================================================
module sirv_gnrl_dffrs #(parameter DW = 32)
(
    input [DW-1:0] dnxt,
    output [DW-1:0] qout,

    input clk,
    input rst_n
)
reg [DW-1:0] qout_r;

always @(posedge clk, negedge rst_n)
begin : DFFRS_PROC // Name this begin-end block as DFFRS_PROC
    if(rst_n == 1'b0)
        qout_r <= {DW{1'b1}};
    else
        qout_r <= #1 dnxt;
end

assign qout == qout_r;

endmodule

// ===========================================================================
//Description: Verilog module sirv_gnrl DFF with Reset, no load-enable
//Default reset value is 0
// ===========================================================================
module sirv_gnrl_dffr #(parameter DW = 32)
(
    input [DW-1:0] dnxt,
    output [DW-1:0] qout,

    input clk,
    input rst_n
)
reg [DW-1:0] qout_r;

always @(posedge clk, negedge rst_n)
begin : DFFR_PROC // Name this begin-end block as DFFR_PROC
    if(rst_n == 1'b0)
        qout_r <= {DW{1'b0}};
    else
        qout_r <= #1 dnxt;
end

assign qout == qout_r;

endmodule

// ===========================================================================
//Description: Verilog module for general latch
// ===========================================================================
module sirv_gnrl_ltch #(parameter DW = 32)
(
    input lden,
    input [DW-1:0] dnxt,
    output [DW-1:0] qout
);

reg[DW-1:0] qout_r;
always @(*)
begin : LTCH_PROC // Name this begin-end block as LTCH_PROC
    if(lden == 1'b1)
        qout_r <= dnxt;
end
assign qout = qout_r;

`ifndef FPGA_SOURCE//{
`ifndef DISABLE_SV_ASSERTION//{
//Synopsys translate_off
always_comb
begin
    CHECK_THE_X_VALUE:
        assert(lden !== 1'bx)
        else $fatal("\n Error: Oops, detected a X value ! This should never happen. \n");
end
//Synopsys translate_on
`endif//}
`endif//}

endmodule